module crud

import os
import mysql

// create user
pub fn create(api_name string) {

}

pub fn read(api_name string) {

}

pub fn update(api_name string) {

}

pub fn delete(api_name string) {
    
}
