module term_control

import os

pub const (
	// All ANSI Colors Here
)

// Gradient Text
pub fn rgb_text() {

}