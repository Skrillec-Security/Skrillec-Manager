module api_server