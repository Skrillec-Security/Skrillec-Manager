module crud

import os
import mysql

// create user
pub fn create(spoof_ip string) {

}

pub fn read(spoof_ip string) {

}

pub fn update(spoof_ip string) {

}

pub fn delete(spoof_ip string) {
    
}
