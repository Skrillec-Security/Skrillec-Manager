module manager

import os

pub fn cmd_handler(cmd string) {

}