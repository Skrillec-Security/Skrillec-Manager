module crud

import os
import mysql

// create user
pub fn create(key string) {

}

pub fn read(key string) {

}

pub fn update(key string) {

}

pub fn delete(key string) {
    
}
